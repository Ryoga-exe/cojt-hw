//-----------------------------------------------------------------------------
// Module : tb_led7_dec
//-----------------------------------------------------------------------------
`timescale 1ns / 1ns

module tb_led7_dec;

  //-----------------------------------------------------------------------------
  //	Internal Signals
  //-----------------------------------------------------------------------------
  logic [3:0] disp_data;  //display data
  logic disp_en;  //display enable
  logic [6:0] segment;  //7segment data active low

  //-----------------------------------------------------------------------------
  //	Parameter Definition
  //-----------------------------------------------------------------------------
  // simulation step
  parameter STEP = 10;

  //-----------------------------------------------------------------------------
  //	Module Call
  //-----------------------------------------------------------------------------
  led7_dec i_led7_dec (
      .disp_data(disp_data),
      .disp_en  (disp_en),
      .segment  (segment)
  );

  //-----------------------------------------------------------------------------
  //	Clock Generate
  //-----------------------------------------------------------------------------

  //-----------------------------------------------------------------------------
  //	Simulation
  //-----------------------------------------------------------------------------
  integer i;

  initial begin
    // set initial value
    disp_data = 4'd0;
    disp_en   = 1'b0;

    // test 1
    disp_en   = 1'b1;
    for (i = 0; i < 16; i = i + 1) begin
      disp_data = i[3:0];
      #STEP;
    end

    repeat (5) #STEP;

    // test 2
    disp_en = 1'b0;
    for (i = 0; i < 15; i = i + 1) begin
      disp_data = i[3:0];
      #STEP;
    end

    repeat (5) #STEP;

    $display("-----------------------------------------\n");
    $display("            Simulation  Finish !!        \n");
    $display("-----------------------------------------\n");
    $finish;
  end

endmodule
