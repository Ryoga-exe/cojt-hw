//-----------------------------------------------------------------------------
// Module : tb_en_gen
//-----------------------------------------------------------------------------
`timescale 1ns/1ns

module tb_en_gen;

//-----------------------------------------------------------------------------
//	Internal Signals
//-----------------------------------------------------------------------------
logic			clk;					// system clk
logic			rst;					// synchronous reset

logic			en_1hz;					// 1Hz enable out
logic			mask_1hz;				// 1Hz blinking out

//-----------------------------------------------------------------------------
//	Parameter Definition
//-----------------------------------------------------------------------------
// CLK = 100MHz : 10ns/T
parameter cycle = 10;

//-----------------------------------------------------------------------------
//	Module Call
//-----------------------------------------------------------------------------
en_gen		i_en_gen(
	.clk		(clk),
	.rst		(rst),
	.en_1hz		(en_1hz),
	.mask_1hz	(mask_1hz) );

//-----------------------------------------------------------------------------
//	Clock Generate
//-----------------------------------------------------------------------------
always begin
	clk = 1'b0;
	#(cycle/2);
	clk = 1'b1;
	#(cycle/2);
end

//-----------------------------------------------------------------------------
//	Simulation
//-----------------------------------------------------------------------------
initial begin
// set initial value
	rst = 1'b0;

// reset in
	TASK_RESET;
	@(posedge clk);

// test of free run count up 
	repeat (159999999) @(posedge clk);

	$display("-----------------------------------------\n");
	$display("            Simulation  Finish !!        \n");
	$display("-----------------------------------------\n");
	$finish;
end

//-----------------------------------------------------------------------------
//	Task Definition
//-----------------------------------------------------------------------------
task TASK_RESET;
	@(posedge clk);
	#(1);
	rst= 1'b1 ;
	repeat(3) @(posedge clk);
	#(1);
	rst = 1'b0;
endtask

endmodule


